`timescale 1ns / 1ps
`default_nettype none

`ifdef SYNTHESIS
`define FPATH(X) `"X`"
`else /* ! SYNTHESIS */
`define FPATH(X) `"../../data/X`"
`endif  /* ! SYNTHESIS */

module image_sprite #(
  parameter WIDTH=256, HEIGHT=256) (
  input wire pixel_clk_in,
  input wire rst_in,
  input wire pop_in, // 0: closed, 1: open 
  input wire [10:0] x_in, hcount_in,
  input wire [9:0]  y_in, vcount_in,
  output logic [7:0] red_out,
  output logic [7:0] green_out,
  output logic [7:0] blue_out
  );
  // open mouth no offset
  // closed mouth +offset

  // calculate rom address
  logic [$clog2(WIDTH*HEIGHT*2+1)-1:0] image_addr;
  logic [$clog2(WIDTH*HEIGHT*2+1)-1:0] sprite_offset;
  assign sprite_offset = pop_in ? 0 : 256*256;
  assign image_addr = (hcount_in - x_in) + ((vcount_in - y_in) * WIDTH) + sprite_offset;

  logic in_sprite, in_sprite_pipelined;
  assign in_sprite = ((hcount_in >= x_in && hcount_in < (x_in + WIDTH)) &&
                      (vcount_in >= y_in && vcount_in < (y_in + HEIGHT)));

  pipeline #(.STAGES(4)) isp(.clk_in(pixel_clk_in), .sig_in(in_sprite), .sig_out(in_sprite_pipelined));
  // Modify the module below to use your BRAMs!
  assign red_out =    in_sprite_pipelined ? palette_out[23:16] : 0;
  assign green_out =  in_sprite_pipelined ? palette_out[15:8] : 0;
  assign blue_out =   in_sprite_pipelined ? palette_out[7:0] : 0;

  logic [23:0] palette_out;
  logic [7:0] image_out;

  xilinx_single_port_ram_read_first #(
    .RAM_WIDTH(8),                       // Specify RAM data width
    .RAM_DEPTH(256*256*2),                     // Specify RAM depth (number of entries)
    .RAM_PERFORMANCE("HIGH_PERFORMANCE"), // Select "HIGH_PERFORMANCE" or "LOW_LATENCY" 
    .INIT_FILE(`FPATH(image2.mem))          // Specify name/location of RAM initialization file if using one (leave blank if not)
  ) image_mem (
    .addra(image_addr),     // Address bus, width determined from RAM_DEPTH
    .dina(0),       // RAM input data, width determined from RAM_WIDTH
    .clka(pixel_clk_in),       // Clock
    .wea(0),         // Write enable
    .ena(1),         // RAM Enable, for additional power savings, disable port when not in use
    .rsta(rst_in),       // Output reset (does not affect memory contents)
    .regcea(1),   // Output register enable
    .douta(image_out)      // RAM output data, width determined from RAM_WIDTH
  );

  xilinx_single_port_ram_read_first #(
    .RAM_WIDTH(8*3),                      // Specify RAM data width
    .RAM_DEPTH(256),                      // Specify RAM depth (number of entries)
    .RAM_PERFORMANCE("HIGH_PERFORMANCE"), // Select "HIGH_PERFORMANCE" or "LOW_LATENCY" 
    .INIT_FILE(`FPATH(palette2.mem))      // Specify name/location of RAM initialization file if using one (leave blank if not)
  ) palette_mem (
    .addra(image_out),     // Address bus, width determined from RAM_DEPTH
    .dina(0),       // RAM input data, width determined from RAM_WIDTH
    .clka(pixel_clk_in),       // Clock
    .wea(0),         // Write enable
    .ena(1),         // RAM Enable, for additional power savings, disable port when not in use
    .rsta(rst_in),       // Output reset (does not affect memory contents)
    .regcea(1),   // Output register enable
    .douta(palette_out)      // RAM output data, width determined from RAM_WIDTH
  );


endmodule






`default_nettype none
